`ifndef DEFINES_VH
`define DEFINES_VH

`define DATA_WIDTH 8
`define ACC_WIDTH 20

`endif
